// gps_connection.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module gps_connection (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

endmodule
